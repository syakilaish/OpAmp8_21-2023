* Created by KLayout

* cell Op8_18_rev1
* pin Out
* pin Bias
* pin Vdd
* pin In+
* pin In1
* pin Vss
.SUBCKT Op8_18_rev1 4 14 16 18 21 25
* net 4 Out
* net 14 Bias
* net 16 Vdd
* net 18 In+
* net 21 In1
* net 25 Vss
* device instance $1 r0 *1 109,44 NMOS
M$1 2 1 25 25 NMOS L=5U W=20U AS=30P AD=30P PS=36U PD=36U
* device instance $3 r0 *1 148,44 NMOS
M$3 4 3 25 25 NMOS L=1U W=100U AS=110P AD=110P PS=132U PD=132U
* device instance $13 m90 *1 138,44 NMOS
M$13 5 5 25 25 NMOS L=1U W=40U AS=50P AD=50P PS=60U PD=60U
* device instance $17 m90 *1 138,62 NMOS
M$17 8 8 5 25 NMOS L=1U W=40U AS=50P AD=50P PS=60U PD=60U
* device instance $21 m90 *1 145.5,103 NMOS
M$21 17 8 3 25 NMOS L=1U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $26 m90 *1 82,44 NMOS
M$26 6 11 25 25 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $27 r0 *1 95.5,44 NMOS
M$27 7 11 25 25 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $28 m90 *1 57,127.5 NMOS
M$28 19 18 13 25 NMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $33 r0 *1 67.5,127.5 NMOS
M$33 20 21 13 25 NMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $38 r0 *1 42,79 NMOS
M$38 13 12 10 25 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $43 m90 *1 32,49 NMOS
M$43 9 1 25 25 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $48 r0 *1 42,49 NMOS
M$48 10 1 25 25 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $53 r0 *1 93.5,69 NMOS
M$53 3 11 7 25 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $58 m90 *1 84,69 NMOS
M$58 11 11 6 25 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $63 m90 *1 32,79 NMOS
M$63 1 12 9 25 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $68 r0 *1 112.5,190.5 PMOS
M$68 8 14 16 16 PMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $69 r0 *1 148.5,165.5 PMOS
M$69 4 17 16 16 PMOS L=1U W=600U AS=660P AD=660P PS=682U PD=682U
* device instance $79 m90 *1 133.5,152.5 PMOS
M$79 2 2 22 16 PMOS L=1U W=80U AS=100P AD=100P PS=110U PD=110U
* device instance $83 m90 *1 136,185.5 PMOS
M$83 22 22 16 16 PMOS L=1U W=80U AS=100P AD=100P PS=110U PD=110U
* device instance $87 m90 *1 119.5,107.5 PMOS
M$87 3 2 17 16 PMOS L=1U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $92 r0 *1 40,161 PMOS
M$92 12 14 24 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $97 r0 *1 41.5,187.5 PMOS
M$97 24 14 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $99 r0 *1 91.5,188 PMOS
M$99 19 14 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $101 r0 *1 71.5,188 PMOS
M$101 20 14 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $103 r0 *1 69,160.5 PMOS
M$103 11 14 20 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $108 m90 *1 30,161 PMOS
M$108 14 14 23 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $113 r0 *1 96,160.5 PMOS
M$113 17 14 19 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $118 m90 *1 28.5,187.5 PMOS
M$118 23 14 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $120 r90 *1 78.5,103.5 HRES
R$120 12 1 17500 HRES
* device instance $123 r270 *1 37.5,103.5 HRES
R$123 25 14 350000 HRES
* device instance $125 m45 *1 164,75.5 CAP
C$125 4 3 1.56e-12 CAP
* device instance $126 r270 *1 164,109.5 CAP
C$126 4 17 1.56e-12 CAP
.ENDS Op8_18_rev1
