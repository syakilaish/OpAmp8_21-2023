* Created by KLayout

* cell TOP
* pin Out
* pin Ibias
* pin Vdd
* pin Vss
.SUBCKT TOP 4 15 16 22
* net 4 Out
* net 15 Ibias
* net 16 Vdd
* net 22 Vss
* device instance $1 r0 *1 109,44 NMOS
M$1 2 1 22 22 NMOS L=5U W=20U AS=30P AD=30P PS=36U PD=36U
* device instance $3 r0 *1 147,44 NMOS
M$3 4 3 22 22 NMOS L=1U W=100U AS=110P AD=110P PS=132U PD=132U
* device instance $13 m90 *1 138,44 NMOS
M$13 5 5 22 22 NMOS L=1U W=40U AS=50P AD=50P PS=60U PD=60U
* device instance $17 m90 *1 138,62 NMOS
M$17 8 8 5 22 NMOS L=1U W=40U AS=50P AD=50P PS=60U PD=60U
* device instance $21 m90 *1 136.5,103.5 NMOS
M$21 14 8 3 22 NMOS L=1U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $26 m90 *1 82,44 NMOS
M$26 6 12 22 22 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $27 r0 *1 95.5,44 NMOS
M$27 7 12 22 22 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $28 r0 *1 42,79 NMOS
M$28 13 11 10 22 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $33 m90 *1 32,49 NMOS
M$33 9 1 22 22 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $38 r0 *1 42,49 NMOS
M$38 10 1 22 22 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $43 r0 *1 93.5,69 NMOS
M$43 3 12 7 22 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $48 m90 *1 84,69 NMOS
M$48 12 12 6 22 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $53 m90 *1 57,130 NMOS
M$53 17 23 13 22 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $58 r0 *1 65,130 NMOS
M$58 18 24 13 22 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $63 m90 *1 32,79 NMOS
M$63 1 11 9 22 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $68 r0 *1 112.5,190.5 PMOS
M$68 8 15 16 16 PMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $69 r0 *1 148.5,165.5 PMOS
M$69 4 14 16 16 PMOS L=1U W=600U AS=660P AD=660P PS=682U PD=682U
* device instance $79 m90 *1 133.5,152.5 PMOS
M$79 2 2 19 16 PMOS L=1U W=80U AS=100P AD=100P PS=110U PD=110U
* device instance $83 m90 *1 136,185.5 PMOS
M$83 19 19 16 16 PMOS L=1U W=80U AS=100P AD=100P PS=110U PD=110U
* device instance $87 m90 *1 109.5,116.5 PMOS
M$87 3 2 14 16 PMOS L=1U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $92 r0 *1 41.5,187.5 PMOS
M$92 21 15 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $94 r0 *1 71.5,188 PMOS
M$94 18 15 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $96 r0 *1 91.5,188 PMOS
M$96 17 15 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $98 r0 *1 40,161 PMOS
M$98 11 15 21 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $103 r0 *1 69,160.5 PMOS
M$103 12 15 18 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $108 r0 *1 96,160.5 PMOS
M$108 14 15 17 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $113 m90 *1 30,161 PMOS
M$113 15 15 20 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $118 m90 *1 28.5,187.5 PMOS
M$118 20 15 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $120 r180 *1 16.5,120.5 HRES
R$120 22 15 350000 HRES
* device instance $124 r90 *1 52,106 HRES
R$124 11 1 17500 HRES
* device instance $125 m45 *1 161.5,75.5 CAP
C$125 4 3 1.56e-12 CAP
* device instance $126 r270 *1 161.5,109.5 CAP
C$126 4 14 1.56e-12 CAP
.ENDS TOP
