* Created by KLayout

* cell Op8_18
* pin Out
* pin Vdd
* pin Bias
* pin Vss
.SUBCKT Op8_18 4 16 19 23
* net 4 Out
* net 16 Vdd
* net 19 Bias
* net 23 Vss
* device instance $1 r0 *1 109,44 NMOS
M$1 2 1 23 23 NMOS L=5U W=20U AS=30P AD=30P PS=36U PD=36U
* device instance $3 r0 *1 147,44 NMOS
M$3 4 3 23 23 NMOS L=1U W=100U AS=110P AD=110P PS=132U PD=132U
* device instance $13 m90 *1 138,44 NMOS
M$13 5 5 23 23 NMOS L=1U W=40U AS=50P AD=50P PS=60U PD=60U
* device instance $17 m90 *1 138,62 NMOS
M$17 8 8 5 23 NMOS L=1U W=40U AS=50P AD=50P PS=60U PD=60U
* device instance $21 m90 *1 141.5,103 NMOS
M$21 15 8 3 23 NMOS L=1U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $26 m90 *1 82,44 NMOS
M$26 6 11 23 23 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $27 r0 *1 95.5,44 NMOS
M$27 7 11 23 23 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $28 m90 *1 55.5,127 NMOS
M$28 17 24 13 23 NMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $33 r0 *1 66.5,127 NMOS
M$33 18 25 13 23 NMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $38 r0 *1 42,79 NMOS
M$38 13 12 10 23 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $43 m90 *1 32,49 NMOS
M$43 9 1 23 23 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $48 r0 *1 42,49 NMOS
M$48 10 1 23 23 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $53 r0 *1 93.5,69 NMOS
M$53 3 11 7 23 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $58 m90 *1 84,69 NMOS
M$58 11 11 6 23 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $63 m90 *1 32,79 NMOS
M$63 1 12 9 23 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $68 r0 *1 112.5,190.5 PMOS
M$68 8 19 16 16 PMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $69 r0 *1 148.5,165.5 PMOS
M$69 4 15 16 16 PMOS L=1U W=600U AS=660P AD=660P PS=682U PD=682U
* device instance $79 m90 *1 133.5,152.5 PMOS
M$79 2 2 20 16 PMOS L=1U W=80U AS=100P AD=100P PS=110U PD=110U
* device instance $83 m90 *1 136,185.5 PMOS
M$83 20 20 16 16 PMOS L=1U W=80U AS=100P AD=100P PS=110U PD=110U
* device instance $87 m90 *1 119.5,107.5 PMOS
M$87 3 2 15 16 PMOS L=1U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $92 r0 *1 41.5,187.5 PMOS
M$92 22 19 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $94 r0 *1 91.5,188 PMOS
M$94 17 19 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $96 r0 *1 71.5,188 PMOS
M$96 18 19 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $98 r0 *1 69,160.5 PMOS
M$98 11 19 18 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $103 r0 *1 40,161 PMOS
M$103 12 19 22 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $108 r0 *1 96,160.5 PMOS
M$108 15 19 17 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $113 m90 *1 30,161 PMOS
M$113 19 19 21 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $118 m90 *1 28.5,187.5 PMOS
M$118 21 19 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $120 r90 *1 78.5,103.5 HRES
R$120 12 1 11666.6666667 HRES
* device instance $123 r270 *1 37.5,101.75 HRES
R$123 23 19 186666.666667 HRES
* device instance $125 m45 *1 161.5,75.5 CAP
C$125 28 3 1.56e-12 CAP
* device instance $126 r270 *1 161.5,109.5 CAP
C$126 29 15 1.56e-12 CAP
.ENDS Op8_18
